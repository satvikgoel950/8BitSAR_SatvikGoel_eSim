// Code created by satvikgoel950@gmail.com
module buff8bit(output [7:0] out, input[7:0]in);
  assign out=in;
endmodule